library verilog;
use verilog.vl_types.all;
entity Enes_Sahin_2018510093_DEUNIAC is
    port(
        V               : out    vl_logic;
        ALU_OPR         : out    vl_logic_vector(2 downto 0);
        out_IR          : out    vl_logic_vector(10 downto 0);
        IR_load         : out    vl_logic;
        T2              : out    vl_logic;
        SC_clear        : out    vl_logic;
        D8              : out    vl_logic;
        T4              : out    vl_logic;
        D10             : out    vl_logic;
        D9              : out    vl_logic;
        T6              : out    vl_logic;
        Q               : out    vl_logic;
        clk             : in     vl_logic;
        D7              : out    vl_logic;
        D11             : out    vl_logic;
        D13             : out    vl_logic;
        T5              : out    vl_logic;
        D12             : out    vl_logic;
        D14             : out    vl_logic;
        T7              : out    vl_logic;
        D15             : out    vl_logic;
        D0              : out    vl_logic;
        D2              : out    vl_logic;
        D1              : out    vl_logic;
        D3              : out    vl_logic;
        D5              : out    vl_logic;
        D4              : out    vl_logic;
        D6              : out    vl_logic;
        out_IM          : out    vl_logic_vector(10 downto 0);
        T0              : out    vl_logic;
        out_PC          : out    vl_logic_vector(4 downto 0);
        PC_count_en     : out    vl_logic;
        T3              : out    vl_logic;
        out_AR          : out    vl_logic_vector(3 downto 0);
        AR_load         : out    vl_logic;
        out_SM          : out    vl_logic_vector(4 downto 0);
        out_SP          : out    vl_logic_vector(3 downto 0);
        R0_out          : out    vl_logic_vector(3 downto 0);
        R0_ld           : out    vl_logic;
        out_BUS         : out    vl_logic_vector(3 downto 0);
        BUS_data_sel    : out    vl_logic;
        out_DM          : out    vl_logic_vector(3 downto 0);
        DM_write        : out    vl_logic;
        DM_read         : out    vl_logic;
        R1_out          : out    vl_logic_vector(3 downto 0);
        R1_ld           : out    vl_logic;
        R2_out          : out    vl_logic_vector(3 downto 0);
        R2_ld           : out    vl_logic;
        InpR_out        : out    vl_logic_vector(3 downto 0);
        input_InpR      : in     vl_logic_vector(3 downto 0);
        out_alu         : out    vl_logic_vector(3 downto 0);
        BUS_sel         : out    vl_logic_vector(1 downto 0);
        T1              : out    vl_logic;
        OUTR_load       : out    vl_logic;
        out_SC          : out    vl_logic_vector(2 downto 0);
        OutpR_out       : out    vl_logic_vector(3 downto 0)
    );
end Enes_Sahin_2018510093_DEUNIAC;
