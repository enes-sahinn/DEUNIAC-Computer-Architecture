library verilog;
use verilog.vl_types.all;
entity Enes_Sahin_2018510093_DEUNIAC_vlg_vec_tst is
end Enes_Sahin_2018510093_DEUNIAC_vlg_vec_tst;
