library verilog;
use verilog.vl_types.all;
entity Enes_Sahin_2018510093_DEUNIAC_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        input_InpR      : in     vl_logic_vector(3 downto 0);
        sampler_tx      : out    vl_logic
    );
end Enes_Sahin_2018510093_DEUNIAC_vlg_sample_tst;
