library verilog;
use verilog.vl_types.all;
entity Enes_Sahin_2018510093_Asgn1_vlg_check_tst is
    port(
        out_alu         : in     vl_logic_vector(3 downto 0);
        overflow        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Enes_Sahin_2018510093_Asgn1_vlg_check_tst;
