library verilog;
use verilog.vl_types.all;
entity Enes_Sahin_2018510093_DEUNIAC_vlg_check_tst is
    port(
        ALU_OPR         : in     vl_logic_vector(2 downto 0);
        AR_load         : in     vl_logic;
        BUS_data_sel    : in     vl_logic;
        BUS_sel         : in     vl_logic_vector(1 downto 0);
        D0              : in     vl_logic;
        D1              : in     vl_logic;
        D2              : in     vl_logic;
        D3              : in     vl_logic;
        D4              : in     vl_logic;
        D5              : in     vl_logic;
        D6              : in     vl_logic;
        D7              : in     vl_logic;
        D8              : in     vl_logic;
        D9              : in     vl_logic;
        D10             : in     vl_logic;
        D11             : in     vl_logic;
        D12             : in     vl_logic;
        D13             : in     vl_logic;
        D14             : in     vl_logic;
        D15             : in     vl_logic;
        DM_read         : in     vl_logic;
        DM_write        : in     vl_logic;
        InpR_out        : in     vl_logic_vector(3 downto 0);
        IR_load         : in     vl_logic;
        out_alu         : in     vl_logic_vector(3 downto 0);
        out_AR          : in     vl_logic_vector(3 downto 0);
        out_BUS         : in     vl_logic_vector(3 downto 0);
        out_DM          : in     vl_logic_vector(3 downto 0);
        out_IM          : in     vl_logic_vector(10 downto 0);
        out_IR          : in     vl_logic_vector(10 downto 0);
        out_PC          : in     vl_logic_vector(4 downto 0);
        out_SC          : in     vl_logic_vector(2 downto 0);
        out_SM          : in     vl_logic_vector(4 downto 0);
        out_SP          : in     vl_logic_vector(3 downto 0);
        OutpR_out       : in     vl_logic_vector(3 downto 0);
        OUTR_load       : in     vl_logic;
        PC_count_en     : in     vl_logic;
        Q               : in     vl_logic;
        R0_ld           : in     vl_logic;
        R0_out          : in     vl_logic_vector(3 downto 0);
        R1_ld           : in     vl_logic;
        R1_out          : in     vl_logic_vector(3 downto 0);
        R2_ld           : in     vl_logic;
        R2_out          : in     vl_logic_vector(3 downto 0);
        SC_clear        : in     vl_logic;
        T0              : in     vl_logic;
        T1              : in     vl_logic;
        T2              : in     vl_logic;
        T3              : in     vl_logic;
        T4              : in     vl_logic;
        T5              : in     vl_logic;
        T6              : in     vl_logic;
        T7              : in     vl_logic;
        V               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Enes_Sahin_2018510093_DEUNIAC_vlg_check_tst;
